library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.aux_package.ALL;

-----------------------------------------
-- Entity Declaration for FIR Filter
-----------------------------------------
entity FIR_Filter is
    Port (
        -- Clock and Reset
        FIRCLK   : in  STD_LOGIC;          -- FIR core clock
        FIFOCLK  : in  STD_LOGIC;          -- FIFO clock
        FIRRST   : in  STD_LOGIC;          -- FIR core reset
        FIFORST  : in  STD_LOGIC;          -- FIFO reset
        
        -- Control signals
        FIRENA   : in  STD_LOGIC;          -- FIR core enable
        FIFOWEN  : in  STD_LOGIC;          -- FIFO write enable
        FIFOREN  : in  STD_LOGIC;          -- FIFO read enable
        
        -- Status signals
        FIFOFULL : out STD_LOGIC;          -- FIFO full status
        FIFOEMPTY: out STD_LOGIC;          -- FIFO empty status
        FIRIFG   : out STD_LOGIC;          -- FIR interrupt flag
        FIRIFG_OUTREADY : out std_logic;   -- NEW: asserts when FIROUT is valid

        -- Data interface
        FIRIN  : in  STD_LOGIC_VECTOR(31 downto 0);   -- FIR input data
        FIROUT : out STD_LOGIC_VECTOR(31 downto 0);   -- FIR output data
        
        -- Coefficient interface
        COEF0 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF1 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF2 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF3 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF4 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF5 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF6 : in STD_LOGIC_VECTOR(7 downto 0);
        COEF7 : in STD_LOGIC_VECTOR(7 downto 0);
        
        -- Memory interface
        Addr     : in STD_LOGIC_VECTOR(11 DOWNTO 0);
        FIRRead  : in STD_LOGIC;
        FIRWrite : in STD_LOGIC;
        
        -- Interrupt control
        FIRIFG_CLR : in STD_LOGIC
    );
end FIR_Filter;

----------------------------------------
-- Architecture Definition
----------------------------------------
architecture Behavioral of FIR_Filter is
    -- Constants
    constant M : integer := 8;  -- Number of filter taps
    constant W : integer := 24; -- Data width
    constant q : integer := 8;  -- Coefficient width
    constant k : integer := 8;  -- FIFO depth parameter
    
    -- FIFO signals
    type fifo_array is array (0 to 2**k-1) of STD_LOGIC_VECTOR(W-1 downto 0);
    signal fifo_memory : fifo_array := (others => (others => '0'));
    signal fifo_wr_ptr : integer range 0 to 2**k-1 := 0;
    signal fifo_rd_ptr : integer range 0 to 2**k-1 := 0;
    signal fifo_count_wr : integer range 0 to 2**k := 0;
    signal fifo_count_rd : integer range 0 to 2**k := 0;
    signal fifo_count    : integer range 0 to 2**k := 0;
    
    -- FIR filter signals
    type delay_line is array (0 to M-1) of STD_LOGIC_VECTOR(W-1 downto 0);
    type coeff_array is array (0 to M-1) of STD_LOGIC_VECTOR(31 downto 0);
    signal x_delay : delay_line := (others => (others => '0'));
    signal coefficients : coeff_array := (others => (others => '0'));
    
    -- Processing signals
    signal x_input : STD_LOGIC_VECTOR(W-1 downto 0);
    signal y_output : STD_LOGIC_VECTOR(31 downto 0);
    signal processing_active : STD_LOGIC := '0';
    
    -- Internal status
    signal fifo_empty_internal : STD_LOGIC;
    signal fifo_full_internal  : STD_LOGIC;
    signal output_valid : std_logic := '0';
    
begin
    ----------------------------------------------------------------
    -- Concurrent assignments 
    ----------------------------------------------------------------
    fifo_empty_internal <= '1' when fifo_count = 0 else '0';
    fifo_full_internal  <= '1' when fifo_count = 2**k-1 else '0';
    
    FIFOEMPTY <= fifo_empty_internal;
    FIFOFULL  <= fifo_full_internal;

    ----------------------------------------------------------------
    -- FIFO write process
    ----------------------------------------------------------------
    process(FIFOCLK, FIFORST)
    begin
        if FIFORST = '1' then
            fifo_wr_ptr   <= 0;
            fifo_count_wr <= 0;
        elsif rising_edge(FIFOCLK) then
            if FIFOWEN = '1' and fifo_count < 2**k-1 then
                fifo_memory(fifo_wr_ptr) <= FIRIN(W-1 downto 0);
                fifo_wr_ptr   <= (fifo_wr_ptr + 1) mod 2**k;
                fifo_count_wr <= fifo_count_wr + 1;
            end if;
        end if;
    end process;

    ----------------------------------------------------------------
    -- FIFO read process (directly uses FIFOREN now)
    ----------------------------------------------------------------
    process(FIRCLK, FIRRST)
    begin
        if FIRRST = '1' then
            fifo_rd_ptr   <= 0;
            x_input       <= (others => '0');
            fifo_count_rd <= 0;
        elsif rising_edge(FIRCLK) then
            if FIFOREN = '1' and fifo_count > 0 then
                x_input       <= fifo_memory(fifo_rd_ptr);
                fifo_rd_ptr   <= (fifo_rd_ptr + 1) mod 2**k;
                fifo_count_rd <= fifo_count_rd + 1;
            end if;
        end if;
    end process;

    ----------------------------------------------------------------
    -- FIFO count combine
    ----------------------------------------------------------------
    fifo_count <= fifo_count_wr - fifo_count_rd;

    ----------------------------------------------------------------
    -- Coefficients
    ----------------------------------------------------------------
    coefficients(0) <= "000000000000000000000000" & COEF0;
    coefficients(1) <= "000000000000000000000000" & COEF1;
    coefficients(2) <= "000000000000000000000000" & COEF2;
    coefficients(3) <= "000000000000000000000000" & COEF3;
    coefficients(4) <= "000000000000000000000000" & COEF4;
    coefficients(5) <= "000000000000000000000000" & COEF5;
    coefficients(6) <= "000000000000000000000000" & COEF6;
    coefficients(7) <= "000000000000000000000000" & COEF7;

    ----------------------------------------------------------------
    -- FIR compute
    ----------------------------------------------------------------
    process(FIRCLK, FIRRST)
        variable temp_sum : signed(55 downto 0);
    begin
        if FIRRST = '1' then
            x_delay          <= (others => (others => '0'));
            y_output         <= (others => '0');
            processing_active <= '0';
        elsif rising_edge(FIRCLK) then
            if FIRENA = '1' then
                -- shift
                for i in M-1 downto 1 loop
                    x_delay(i) <= x_delay(i-1);
                end loop;
                x_delay(0) <= x_input;

                -- MAC
                temp_sum := (others => '0');
                for i in 0 to M-1 loop
                    temp_sum := temp_sum + signed(x_delay(i)) * signed(coefficients(i));
                end loop;

                y_output <= std_logic_vector(temp_sum(55 downto 24));
                processing_active <= '1';
            else
                processing_active <= '0';
            end if;
        end if;
    end process;

    ----------------------------------------------------------------
    -- Output valid flag
    ----------------------------------------------------------------
    process(FIRCLK, FIRRST)
    begin
        if FIRRST = '1' then
            output_valid <= '0';
        elsif rising_edge(FIRCLK) then
            if FIRENA = '1' then
                output_valid <= '1';
            else
                output_valid <= '0';
            end if;
        end if;
    end process;

    ----------------------------------------------------------------
    -- Outputs
    ----------------------------------------------------------------
    FIROUT <= "00000000" & y_output(23 downto 0);

    FIRIFG <= '0' when FIRIFG_CLR = '1' else output_valid;
    FIRIFG_OUTREADY <= output_valid;

end Behavioral;
