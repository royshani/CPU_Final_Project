
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE work.aux_package.ALL;
-----------------------------------------
-- Entity Declaration for MCU
-----------------------------------------
ENTITY MCU IS
	GENERIC(MemWidth	: INTEGER := 10;
			SIM 		: BOOLEAN := FALSE;

			CtrlBusSize	: integer := 8;
			AddrBusSize	: integer := 32;
			DataBusSize	: integer := 32;
			IrqSize		: integer := 8;
			RegSize		: integer := 8
			);
	PORT( 
			reset, clock, ena	: IN	STD_LOGIC;
			HEX0, HEX1, HEX2	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX3, HEX4, HEX5	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0);
			LEDR				: OUT	STD_LOGIC_VECTOR(7 DOWNTO 0);
			Switches			: IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
			BTOUT				: OUT   STD_LOGIC;
			KEY1, KEY2, KEY3	: IN	STD_LOGIC);
END MCU;
----------------------------------------
-- Architecture Definition
----------------------------------------
ARCHITECTURE structure OF MCU IS
	SIGNAL resetSim		: STD_LOGIC;
	SIGNAL enaSim		: STD_LOGIC;

	SIGNAL PC			:	STD_LOGIC_VECTOR(9 DOWNTO 0);
	
	-- CHIP SELECT SIGNALS --
	SIGNAL CS_LEDR, CS_SW, CS_KEY		: STD_LOGIC;
	SIGNAL CS_HEX0, CS_HEX1, CS_HEX2	: STD_LOGIC;
	SIGNAL CS_HEX3, CS_HEX4, CS_HEX5, pll_out	: STD_LOGIC;
	SIGNAL CS_FIR		: STD_LOGIC;
	
	
	-- GPIO SIGNALS -- 
	SIGNAL MemReadBus	: 	STD_LOGIC;
	SIGNAL MemWriteBus	:	STD_LOGIC;
	SIGNAL ControlBus	: 	STD_LOGIC_VECTOR(CtrlBusSize-1 DOWNTO 0);
	SIGNAL AddressBus	: 	STD_LOGIC_VECTOR(AddrBusSize-1 DOWNTO 0);
	SIGNAL DataBus		: 	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0);
	
	-- BASIC TIMER --
	SIGNAL BTCTL        : STD_LOGIC_VECTOR(CtrlBusSize-1 DOWNTO 0);
	SIGNAL BTIP         : STD_LOGIC_VECTOR(1 DOWNTO 0); 		-- 2-bit prescaler select (BTCTL(1 downto 0))
	SIGNAL BTCLR        : STD_LOGIC; 							-- Basic Timer Clear strobe (BTCTL(2))
	SIGNAL BTCNT        : STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0);
	SIGNAL BTCCR0       : STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0);
	SIGNAL BTCCR1       : STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0);
	SIGNAL BTIFG        : STD_LOGIC;

	-- FIR Filter signals
	SIGNAL FIRCTL		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL FIRIN		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL FIROUT		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL COEF3_0		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL COEF7_4		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL FIRIFG		:	STD_LOGIC := '0';
	SIGNAL FIRIFG_OUTREADY : STD_LOGIC := '0';  -- NEW: Output ready signal
	SIGNAL FIFOFULL		:	STD_LOGIC := '0';
	SIGNAL FIFOEMPTY	:	STD_LOGIC := '1';
	
	-- FIR Control signals extracted from FIRCTL
	SIGNAL FIRENA		:	STD_LOGIC := '0';  -- FIR core enable (bit 0)
	SIGNAL FIRRST		:	STD_LOGIC := '0';  -- FIR core reset (bit 1)
	SIGNAL FIFOEMPTY_status : STD_LOGIC := '1'; -- FIFO empty status (bit 2, read-only)
	SIGNAL FIFOFULL_status  : STD_LOGIC := '0'; -- FIFO full status (bit 3, read-only)
	SIGNAL FIFORST		:	STD_LOGIC := '0';  -- FIFO reset (bit 4)
	SIGNAL FIFOWEN		:	STD_LOGIC := '0';  -- FIFO write enable (bit 5)
	
	-- DIVIDER signals (commented out to avoid GPIO conflicts with FIR)
	-- SIGNAL DIVIDEND		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	-- SIGNAL DIVISOR		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	-- SIGNAL QUOTIENT		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	-- SIGNAL RESIDUE		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	-- SIGNAL final_QUOTIENT		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	-- SIGNAL final_RESIDUE		:	STD_LOGIC_VECTOR(DataBusSize-1 DOWNTO 0) := (OTHERS => '0');
	-- SIGNAL DIVIFG		:	STD_LOGIC := '0';
	-- SIGNAL DIVENA		:	STD_LOGIC  := '0';
	
	-- INTERRUPT MODULE --
	SIGNAL IntrEn		:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL IFG			:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TypeReg		:	STD_LOGIC_VECTOR(RegSize-1 DOWNTO 0);
	SIGNAL IntrSrc		:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL IRQ_OUT		:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL INTR			:	STD_LOGIC;
	SIGNAL INTA			:	STD_LOGIC;  
	SIGNAL GIE			:	STD_LOGIC;
	SIGNAL INTR_Active	:	STD_LOGIC;
	SIGNAL CLR_IRQ		:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL FIRIFG_CLR	:	STD_LOGIC;
	
	
BEGIN	

	-------------------------- FPGA or ModelSim -----------------------
	resetSim 	<= reset WHEN SIM ELSE not reset;


	
	CPU: MIPS
		GENERIC MAP(
					MemWidth	=> MemWidth,
					SIM 		=> SIM)
		PORT MAP(
					reset		=> resetSim,
					clock		=> pll_out,
					ena			=> ena,
					PC			=> PC,
					ControlBus	=> ControlBus,
					MemReadBus	=> MemReadBus,
					MemWriteBus	=> MemWriteBus,
					AddressBus	=> AddressBus,
					GIE			=> GIE,
					INTR		=> INTR,
					INTA		=> INTA,
					INTR_Active	=> INTR_Active,
					CLR_IRQ		=> CLR_IRQ,
					DataBus		=> DataBus,
					IFG			=> IFG,
					IntrEn      => IntrEn
		);
		
	
	OAD : 	OptAddrDecoder
	PORT MAP(	reset		=> resetSim,
				AddressBus	=> AddressBus(11 DOWNTO 0),
				CS_LEDR		=> CS_LEDR,
				CS_SW		=> CS_SW,
				CS_KEY		=> CS_KEY,
				CS_HEX0		=> CS_HEX0,
				CS_HEX1		=> CS_HEX1,
				CS_HEX2		=> CS_HEX2,
				CS_HEX3		=> CS_HEX3,
				CS_HEX4		=> CS_HEX4,
				CS_HEX5		=> CS_HEX5,
				CS_FIR		=> CS_FIR
				);
		
	
	IO_interface: GPIO
		PORT MAP(
			INTA		=> INTA,
			MemReadBus	=> MemReadBus,
			clock		=> pll_out,
			reset		=> resetSim,
			MemWriteBus	=> MemWriteBus,
			AddressBus	=> AddressBus,
			DataBus		=> DataBus,
			HEX0		=> HEX0,
			HEX1		=> HEX1,
			HEX2		=> HEX2,
			HEX3		=> HEX3,
			HEX4		=> HEX4,
			HEX5		=> HEX5,
			LEDR		=> LEDR,
			Switches	=> Switches,
			CS_LEDR		=> CS_LEDR,
			CS_SW		=> CS_SW,
			CS_HEX0		=> CS_HEX0,
			CS_HEX1		=> CS_HEX1,
			CS_HEX2		=> CS_HEX2,
			CS_HEX3		=> CS_HEX3,
			CS_HEX4		=> CS_HEX4,
			CS_HEX5		=> CS_HEX5
		);

	-- Extract FIR control signals from FIRCTL
	FIRENA <= FIRCTL(0);           -- FIR core enable
	FIRRST <= FIRCTL(1);           -- FIR core reset
	FIFOEMPTY_status <= FIFOEMPTY; -- FIFO empty status (read-only)
	FIFOFULL_status <= FIFOFULL;   -- FIFO full status (read-only)
	FIFORST <= FIRCTL(4);          -- FIFO reset
	FIFOWEN <= FIRCTL(5);          -- FIFO write enable
	
	-- FIR register write process
	PROCESS(pll_out)
	BEGIN
		if (falling_edge(pll_out)) then
			-- Basic Timer registers
			if(AddressBus(11 DOWNTO 0) = X"81C" AND MemWriteBus = '1') then
				BTCTL <= ControlBus;
			END IF;
			
			if(AddressBus(11 DOWNTO 0) = X"824" AND MemWriteBus = '1') then
				BTCCR0 <= DataBus;
			END IF;
			
			if(AddressBus(11 DOWNTO 0) = X"828" AND MemWriteBus = '1') then
				BTCCR1 <= DataBus;
			END IF;
			
			-- FIR registers (handled by FIR component when CS_FIR is active)
			if(CS_FIR = '1' AND MemWriteBus = '1') then
				case AddressBus(11 DOWNTO 0) is
					when X"82C" => FIRCTL <= DataBus;
					when X"830" => FIRIN <= DataBus;
					-- when X"834" => FIROUT <= DataBus;
					when X"838" => COEF3_0 <= DataBus;
					when X"83C" => COEF7_4 <= DataBus;
					when others => null;
				end case;
			end if;
			
			-- DIVIDER registers (commented out to avoid GPIO conflicts)
			-- if(AddressBus(11 DOWNTO 0) = X"82C" AND MemWriteBus = '1') then
			-- 	DIVIDEND <= DataBus;
			-- END IF;
			
			-- if(AddressBus(11 DOWNTO 0) = X"830" AND MemWriteBus = '1') then
			-- 	DIVISOR <= DataBus;
			-- 	DIVENA <= '1';
			-- END IF;
			
			-- if(DIVIFG = '1') then
			-- 	DIVENA <= '0';
			-- 	final_QUOTIENT <= QUOTIENT;
			-- 	final_RESIDUE <= RESIDUE;
			-- END IF;
		END IF;
	END PROCESS;
	
	----
	BTCNT	<= DataBus		WHEN (AddressBus(11 DOWNTO 0) = X"820" AND MemWriteBus = '1') ELSE
			   (OTHERS => 'Z');	-- INPUT

			 
			 
	DataBus <= FIROUT WHEN (AddressBus(11 DOWNTO 0) = X"834" AND MemReadBus = '1')  ELSE
			   -- DIVIDER outputs (commented out to avoid GPIO conflicts)
			   -- final_QUOTIENT WHEN (AddressBus(11 DOWNTO 0) = X"834" AND MemReadBus = '1')  ELSE
			   -- final_RESIDUE WHEN  (AddressBus(11 DOWNTO 0) = X"838" AND MemReadBus = '1')  ELSE
			   "000000000000000000000000" & Switches		WHEN  (AddressBus(11 DOWNTO 0) = X"810" AND MemReadBus = '1')  ELSE
			   "000000000000000000000000"  & IFG WHEN (AddressBus(11 DOWNTO 0) = X"841" AND MemReadBus = '1')  ELSE
			   "000000000000000000000000"  & IntrEn WHEN (AddressBus(11 DOWNTO 0) = X"840" AND MemReadBus = '1')  ELSE
			   BTCNT WHEN (AddressBus(11 DOWNTO 0) = X"820" AND MemReadBus = '1')  ELSE
			   (OTHERS => 'Z');


	-- FIR Filter component
	FIR_acc: FIR_Filter
		Port MAP(
			-- Clock and Reset
			FIRCLK => pll_out,          -- FIR core clock
			FIFOCLK => pll_out,         -- FIFO clock (using same clock for simplicity)
			FIRRST => FIRRST,           -- FIR core reset
			FIFORST => FIFORST,         -- FIFO reset
			
			-- Control signals
			FIRENA => FIRENA,           -- FIR core enable
			FIFOWEN => FIFOWEN,         -- FIFO write enable
			FIFOREN => '1',             -- FIFO read enable (always enabled when processing)
			
			-- Status signals
			FIFOFULL => FIFOFULL,       -- FIFO full status
			FIFOEMPTY => FIFOEMPTY,     -- FIFO empty status
			FIRIFG => FIRIFG,           -- FIR interrupt flag
			FIRIFG_OUTREADY => FIRIFG_OUTREADY, -- NEW: asserts when FIROUT is valid

			-- Data interface
			FIRIN => FIRIN,             -- FIR input data
			FIROUT => FIROUT,           -- FIR output data
			
			-- Coefficient interface
			COEF0 => COEF3_0(7 downto 0),    -- Coefficient 0
			COEF1 => COEF3_0(15 downto 8),   -- Coefficient 1
			COEF2 => COEF3_0(23 downto 16),  -- Coefficient 2
			COEF3 => COEF3_0(31 downto 24),  -- Coefficient 3
			COEF4 => COEF7_4(7 downto 0),    -- Coefficient 4
			COEF5 => COEF7_4(15 downto 8),   -- Coefficient 5
			COEF6 => COEF7_4(23 downto 16),  -- Coefficient 6
			COEF7 => COEF7_4(31 downto 24),  -- Coefficient 7
			
			-- Memory interface
			Addr => AddressBus(11 DOWNTO 0),
			FIRRead => MemReadBus,
			FIRWrite => MemWriteBus,
			
			-- Interrupt control
			FIRIFG_CLR => FIRIFG_CLR    -- Clear FIR interrupt flag
		);

	-- DIVIDER component (commented out to avoid GPIO conflicts)
	-- div_acc: Divider
	-- 	Port MAP(
	-- 		clk => pll_out,          -- Clock signal
	-- 		
	-- 		Addr	=> AddressBus(11 DOWNTO 0),
	-- 		DIVRead	=> MemReadBus,
	-- 		
	-- 		reset => resetSim,       -- Asynchronous reset signal
	-- 		ena  => DIVENA,        -- Start signal to begin the division
	-- 		dividend => DIVIDEND, -- Input for dividend (32-bit)
	-- 		divisor => DIVISOR, -- Input for divisor (32-bit)
	-- 		quotient_OUT => QUOTIENT, -- Output for quotient (32-bit)
	-- 		remainder_OUT => RESIDUE, -- Output for remainder (32-bit)
	-- 		DIVIFG => DIVIFG         -- Indicates an overflow condition
	-- 	);
	
	
	Basic_Timer: BTIMER
		PORT MAP(
			Addr	=> AddressBus(11 DOWNTO 0),
			BTRead	=> MemReadBus,
			BTWrite	=> MemWriteBus,
			MCLK	=> pll_out,
			reset	=> resetSim,
			BTCTL	=> BTCTL,
			BTCCR0	=> BTCCR0,
			BTCCR1	=> BTCCR1,
			BTCNT_io=> BTCNT,
			IRQ_OUT => IRQ_OUT(2),
			BTIFG	=> BTIFG,
			BTOUT	=> BTOUT
		);
		
		
	
	IntrSrc	<=  FIRIFG_OUTREADY  & FIFOEMPTY & (NOT KEY3) & (NOT KEY2) & (NOT KEY1) & BTIFG & '0' & '0';
	Intr_Controller: INTERRUPT
		GENERIC MAP(
			DataBusSize	=> DataBusSize,
			AddrBusSize	=> AddrBusSize,
			IrqSize		=> IrqSize,
			RegSize 	=> RegSize
		)
		PORT MAP(
			reset		=> resetSim,
		    clock		=> pll_out,
		    MemReadBus	=> MemReadBus,
		    MemWriteBus	=> MemWriteBus,
		    AddressBus	=> AddressBus,
		    DataBus		=> DataBus,
		    IntrSrc		=> IntrSrc,
		    ChipSelect	=> '0',
		    INTR		=> INTR,
		    INTA		=> INTA,
			IRQ_OUT		=> IRQ_OUT,
			INTR_Active	=> INTR_Active,
			CLR_IRQ_OUT	=> CLR_IRQ,
		    GIE			=> GIE,
			IFG 		=> IFG,
			IntrEn		=> IntrEn,
			FIRIFG_CLR	=> FIRIFG_CLR
		);
		
		 m1: PLL port map(
	     inclk0 => clock,
		  c0 => pll_out
	   );

	   
	
END structure;